`timescale 1ns/1ps
/*
    A scratchpad memory is a small fast directly accessed RAM used for temporary storage. 
    It is unlike the cache memory where the data is fetched and maintained
    Users directly hardcode values into this memories
*/
module scratchpad(
    
);


endmodule